//interface code 
interface fa_intf;
  logic a,b,s,cin,s,cout;
endinterface
