module test_write;
	initial begin 
	$write("Hello ");
	$write("Amit here.");
	end
endmodule