////test code for the module hello program 
/* module test;
	reg [16*8:0]a;
	
	initial begin 
		a = "Hello World";
		$display("%s, is the string.",a);
	end
endmodule */

/
