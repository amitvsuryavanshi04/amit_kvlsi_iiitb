//code for interface 
interface prio_enco_intf;
  logic [3:0]i;
  logic [1:0]d;
endinterface