module test_monitor;
	initial begin	
		$monitor("Hello");
		$monitor("Amit");
		$monitor("123");
	end
endmodule