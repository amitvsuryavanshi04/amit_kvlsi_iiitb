// Code your design here
module fa(input a,b,cin,output s,cout);
  assign {cout,s} = a+b+cin;
endmodule 
