//binary to gray conversion
interface b2g_intf;
  logic [3:0]bit_in;
  logic [3:0]gray_out;
endinterface