module test;
	initial begin
		$display("Hello");
		$display("Amit Here.");
	end
endmodule