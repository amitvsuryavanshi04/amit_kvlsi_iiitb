// Code your design here
module pattern_numbers_left #(parameter N = 10);  // N is the number of rows
  integer i, j;

  initial begin
    for (i = 1; i <= N; i = i + 1) begin
      for (j = 1; j <= i; j = j + 1) begin
        $write("%0d ", j);
      end
      $display();
    end
  end
endmodule
