//interface 
interface tff_if;
  logic clk, rst;
  logic t;
  logic q;
endinterface